module data_width_converter (
    input clk,
    input resetn,

    input [7:0] data_in,
    input valid_in,
    output ready_in,

    output [23:0] data_out,
    output valid_out,
    input ready_out

);
    
    
endmodule